library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.CPU_library.all;

entity ControlUnit_tb is
end ControlUnit_tb;

architecture Testbench of ControlUnit_tb is

	signal finish_flag		: std_logic := '0';
	constant clk_period		: time := 100 ps;

	component ControlUnit is
	
		port(	
				OpCode		: in std_logic_vector(3 downto 0);
				CLK			: in std_logic;
				Reset			: in std_logic;
				MemtoReg 	: out std_logic;
				GPRF_wr		: out std_logic;
				IR_write 	: out std_logic;
				Mem_wr		: out std_logic;
				Rs2_select	: out std_logic;
				PC_Wcond		: out std_logic;
				Mem_read		: out std_logic;
				PC_write 	: out std_logic;
				PC_source	: out std_logic;
				ALU_op		: out std_logic_vector(3 downto 0);
				ALU_src1		: out std_logic;
				ALU_src2		: out std_logic_vector(1 downto 0);
				Jmp_enable	: out std_logic; 
				IorD			: out std_logic; 
				Cu_state 	: out std_logic_vector(3 downto 0)
		);

	end component;

	signal   OpCode		: std_logic_vector(3 downto 0);
	signal	CLK			: std_logic;
	signal	Reset			: std_logic;
	signal	MemtoReg 	: std_logic;
	signal	GPRF_wr		: std_logic;
	signal	IR_write 	: std_logic;
	signal	Mem_wr		: std_logic;
	signal	Rs2_select	: std_logic;
	signal	PC_Wcond		: std_logic;
	signal	Mem_read		: std_logic;
	signal	PC_write 	: std_logic;
	signal	PC_source	: std_logic;
	signal	ALU_op		: std_logic_vector(3 downto 0);
	signal	ALU_src1		: std_logic;
	signal	ALU_src2		: std_logic_vector(1 downto 0);
	signal	Jmp_enable	: std_logic; 
	signal	IorD			: std_logic; 
	signal	Cu_state 	: std_logic_vector(3 downto 0);
	
	constant TOTAL_CASE	: integer := 10;
	
	type array4bit is array (TOTAL_CASE downto 0) of std_logic_vector(3 downto 0);
	type array2bit is array (TOTAL_CASE downto 0) of std_logic_vector(1 downto 0);
	type array1bit is array (TOTAL_CASE downto 0) of std_logic;
	
	type array2D is array (0 to 15, 0 to 3) of std_logic_vector(3 downto 0); -- 16 opcode and max. 4 states of each 
	constant OpCodeSteps : array2D := (	("0001","0010","0111","1000"), ("0001","0010","0111","1000"), 
													("0001","0010","0111","1000"), ("0001","0010","0111","1000"), 
													("0001","0010","0111","1000"), ("0001","0010","0111","1000"), 
													("0001","0010","0111","1000"), ("0001","0010","0111","1000"),
													("0001","0010","0111","1000"), ("0001","0010","0110","1000"),
													("0001","0010","0110","1111"), ("0001","0010","0011","1111"),
													("0001","0010","1111","1111"), ("0001","0010","0100","1111"),
													("0001","0010","0101","1111"), ("0001","0010","0111","1000"));
													
	type array1D is array (0 to 8) of std_logic_vector(17 downto 0); --control signals total of 18 bit
	constant stateSignals : array1D := ("000000000000000000", "001000110000010100",
													"0000U0000000011000", "000000011000000000",
													"000011001011000010", "000010001011000010",
													"000U00U00000000001", "000000000UUUU0U000",
													"U10000000000000000");

	signal check_enable : std_logic := '0'; -- Check process should perform only when one of the 16 OpCodes occur.
	signal state_signal : integer range 0 to 100 := 1;

	signal 	instruction : STRING (1 TO 7);

	
begin

	UUT: ControlUnit port map(OpCode, CLK, Reset, MemtoReg, GPRF_wr, IR_write, Mem_wr, Rs2_select, PC_Wcond, Mem_read,
										PC_write, PC_source, ALU_op, ALU_src1, ALU_src2, Jmp_enable, IorD, Cu_state) ;
										
										
	Clock: process
	begin
	
		CLK <= '0';
		wait for clk_period/2;
		CLK <= '1';
		wait for clk_period/2;
		
		if finish_flag = '1' then
			wait;
		
		end if; 
	
	end process;
	
	Check: process(CLK, check_enable)
	
		variable state			: integer range 0 to 100 := 1;
		variable OpCodeInt	: integer range 0 to 15 := 0;
		
		variable	MemtoReg_t 		: std_logic;
		variable	GPRF_wr_t		: std_logic;
		variable	IR_write_t 		: std_logic;
		variable	Mem_wr_t			: std_logic;
		variable	Rs2_select_t	: std_logic;
		variable	PC_Wcond_t		: std_logic;
		variable	Mem_read_t		: std_logic;
		variable	PC_write_t 		: std_logic;
		variable	PC_source_t		: std_logic;
		variable	ALU_op_t			: std_logic_vector(3 downto 0);
		variable	ALU_src1_t		: std_logic;
		variable	ALU_src2_t		: std_logic_vector(1 downto 0);
		variable	Jmp_enable_t	: std_logic; 
		variable	IorD_t			: std_logic; 
		
		variable state_temp		: std_logic_vector(17 downto 0);
	
	begin
	
		if falling_edge(CLK) and check_enable = '1' then
			if Cu_state = "0001" then
				state := 0;
				
			else 
				state := state + 1;
				
			end if;
			
			state_signal <= state;
			
			OpCodeInt := to_integer(unsigned(OpCode));
			
			assert Cu_state = OpCodeSteps(OpCodeInt,state)
			report "There is error in OpCode "& integer'image(OpCodeInt) &" and state "& integer'image(state)&" !"
			severity error;
			
			state_temp := stateSignals(to_integer(unsigned(Cu_state)));
			
			MemtoReg_t 		:= state_temp(17);
			GPRF_wr_t 		:= state_temp(16);
			IR_write_t 		:= state_temp(15);
			Mem_wr_t 		:= state_temp(14);
			Rs2_select_t 	:= state_temp(13);
			PC_Wcond_t 		:= state_temp(12);
			Mem_read_t 		:= state_temp(11);
			PC_write_t 		:= state_temp(10);
			PC_source_t 	:= state_temp(9);
			ALU_op_t 		:= state_temp(8 downto 5);
			ALU_src1_t 		:= state_temp(4);
			ALU_src2_t 		:= state_temp(3 downto 2);
			Jmp_enable_t 	:= state_temp(1);
			IorD_t 			:= state_temp(0);
			
		
			case Cu_state is
				
				when "0010" => 
					if OpCode = JZ OR OpCode = JNZ then
						Rs2_select_t := '1';
					else
						Rs2_select_t := '0';
					end if;

				when "0110" => 
					if OpCode = STORE then
						Mem_wr_t := '1';
					else
						Mem_wr_t := '0';
					end if;

					if OpCode = LOAD then
						Mem_read_t := '1';
					else
						Mem_read_t := '0';
					end if;
					
				when "0111" => 

					if OpCode = ADD then
						ALU_op_t := ALU_ADD;
					elsif OpCode = SUBx then
						ALU_op_t := ALU_SUB;
					elsif OpCode = ANDx then
						ALU_op_t := ALU_AND;
					elsif OpCode = ORx then
						ALU_op_t := ALU_OR;
					elsif OpCode = NOTx then
						ALU_op_t := ALU_NOT;
					elsif OpCode = XORx then
						ALU_op_t := ALU_XOR;
					elsif OpCode = CMP then
						ALU_op_t := ALU_CMP;
					elsif OpCode = SHL then
						ALU_op_t := ALU_SHL;
					elsif OpCode = SHR then
						ALU_op_t := ALU_SHR;
					elsif OpCode = LOADI then
						ALU_op_t := ALU_SEL_SRC2;
					end if;

					if OpCode = LOADI then
						ALU_src2_t := "10";
					else
						ALU_src2_t := "00";
					end if;
			
					
				when "1000" => 
					if OpCode = LOAD then
						MemtoReg_t := '1';
					else
						MemtoReg_t := '0';
					end if;
					
				when others => OpCodeInt := to_integer(unsigned(OpCode));
			
			end case;
			
			assert MemtoReg_t = MemtoReg AND GPRF_wr_t = GPRF_wr AND IR_write_t = IR_write AND
					 Mem_wr_t = Mem_wr AND Rs2_select_t = Rs2_select AND PC_Wcond_t = PC_Wcond AND
					 Mem_read_t = Mem_read AND PC_write_t = PC_write AND PC_source_t = PC_source AND
					 ALU_op_t = ALU_op AND ALU_src1_t = ALU_src1 AND ALU_src2_t = ALU_src2 AND
					 Jmp_enable_t = Jmp_enable AND IorD_t = IorD
					 
			report "Errors found in control signals!"
			severity error;
		
		end if;
		
		
	
	end process;
	
	Stimulus: process
	
		variable case_num : integer range 0 to 100 := 1;
	
	begin
	
		Reset <= '1';
		wait for clk_period;
		Reset <= '0';
		wait until Cu_state = "0001";
		
		check_enable <= '1';
		--OpCode <= std_logic_vector(to_unsigned(0,OpCode'length));
		--wait until Cu_state = "0001"; -- Wait until FETCH state.
		for i in 0 to 7 loop --Half of the opcodes
			
			--All opcodes will eventually lead to FETCH state. We need to observe that!
			OpCode <= std_logic_vector(to_unsigned(i,OpCode'length));
			wait until Cu_state = "0001"; -- Wait until FETCH state.
		
		end loop;
		check_enable <= '0';
		
		Reset <= '1';
		wait for clk_period;
		Reset <= '0';
		wait until Cu_state = "0001";
		
		check_enable <= '1';
		for i in 8 to 15 loop --Other half of the opcodes
		
			--All opcodes will eventually lead to FETCH state. We need to observe that!
			OpCode <= std_logic_vector(to_unsigned(i,OpCode'length));
			wait until Cu_state = "0001"; -- Wait until FETCH state.
		
		end loop;
		check_enable <= '0';
		
		finish_flag <= '1';
		wait;
		
	end process;

	IDecoder : PROCESS (OpCode)
	BEGIN
		CASE OpCode IS
			WHEN ADD => 
				instruction <= "ADD    ";
			WHEN SUBx => 
				instruction <= "SUB    ";
			WHEN ANDx => 
				instruction <= "AND    ";
			WHEN ORx => 
				instruction <= "OR     ";
			WHEN NOTx => 
				instruction <= "NOT    ";
			WHEN XORx => 
				instruction <= "XOR    ";
			WHEN CMP => 
				instruction <= "CMP    ";
			WHEN SHL => 
				instruction <= "SHL    ";
			WHEN SHR => 
				instruction <= "SHR    ";
			WHEN LOAD => 
				instruction <= "LOAD   ";
			WHEN STORE => 
				instruction <= "STORE  ";
			WHEN JUMP => 
				instruction <= "JUMP   ";
			WHEN NOP => 
				instruction <= "NOP    ";
			WHEN JZ => 
				instruction <= "JZ     ";
			WHEN JNZ => 
				instruction <= "JNZ    ";
			WHEN LOADI => 
				instruction <= "LOADI  ";			
			WHEN OTHERS => instruction <= "       ";
		END CASE;
	END PROCESS;



end Testbench;